Här är en mening.
Här är en till.