acomp
advcl
advmod
amod
appos
aux
auxpass
cc
ccomp
complm
conj
cop
csubj
csubjpass
dep
det
dobj
expl
infmod
mark
neg
nn
nsubj
nsubjpass
null
num
number
partmod
pcomp
pobj
poss
possessive
preconj
predet
prep
prt
punct
purpcl
quantmod
rcmod
tmod
xcomp
